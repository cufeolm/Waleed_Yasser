`include "add.svh"
`include "add_imm.svh"
`include "and.svh"
`include "and_comp.svh"
`include "and_imm.svh"
`include "and_imm_comp.svh"
`include "xor.svh"
`include "xor_imm.svh"
`include "xor_comp.svh"
`include "xor_imm_comp.svh"
`include "or.svh"
`include "or_imm.svh"
`include "or_comp.svh"
`include "or_imm_comp.svh"
`include "sll.svh"
`include "srl.svh"
`include "sra.svh"

