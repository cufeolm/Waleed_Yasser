`include "GUVM_sequence.sv"
`include "child_sequence.sv"
`include "python_sequence.sv"
`include"add_seq.sv"
`include"bie_seq.sv"
`include"subcc_seq.sv"
