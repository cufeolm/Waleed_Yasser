function void verify_bvsf(GUVM_sequence_item cmd_trans,GUVM_result_transaction res_trans,GUVM_history_transaction hist_trans);
	
	if (cmd_trans.SOM == SB_HISTORY_MODE)
	begin	

		
    end
    
    else if (cmd_trans.SOM == SB_VERIFICATION_MODE)
    begin

	end

endfunction